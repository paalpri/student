paalpri@paalpri.8534:1480330845